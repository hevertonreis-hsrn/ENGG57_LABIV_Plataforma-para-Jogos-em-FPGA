module InstructionMemory (
    input clk,
    //input wire [31:0] address,    // Endereco fornecido pelo PC
    input wire [7:0] address,    // Endereco fornecido pelo PC
    output reg [31:0] instruction // Instrucao de 32 bits lida
);

    // Memoria de instrucoes (256 palavras de 32 bits cada)
    reg [31:0] memory [0:255];

    // Inicialização da memoria com instrucoes (opcional)
    initial begin
        // Carregar algumas instrucoes de exemplo
        memory[0] = 32'b000000_00000_00010_0000000000000001; // LW_1 $2, 1($0)
        memory[1] = 32'b000001_00010_00011_0000000000000000; // LW_2 $3, ($2)
        memory[2] = 32'b000010_00000_00101_0000000000001000; // LW_3 $5, 8
        memory[3] = 32'b000011_00101_00011_0000000000000010; // SW_1 $3, 2($5)
        memory[4] = 32'b000100_00101_00010_0000000000000000; // SW_2 $2, ($5)
        memory[5] = 32'b000101_00011_00100_0000000000000000; // MOV  $4, $3
        memory[6] = 32'b000010_00000_00110_0000000000001010; // LW_3 $6, 10
        memory[7] = 32'b000110_00100_00110_0000000000000000; // ADD  $6, $4
        memory[8] = 32'b000010_00000_00111_0000000000000101; // LW_3 $7, 5
        memory[9] = 32'b000111_00110_00111_0000000000000000; // SUB  $7, $6
        memory[10] = 32'b000010_00000_01000_0000000000000111; // LW_3 $8, 7
        memory[11] = 32'b000010_00000_01001_0000000000001100; // LW_3 $9, 12
        memory[12] = 32'b001000_01000_01001_0000000000000000; // MUL  $9, $8
        memory[13] = 32'b000010_00000_01010_0000000000101100; // LW_3 $10, 44
        memory[14] = 32'b000010_00000_01011_0000000000000010; // LW_3 $11, 2
        memory[15] = 32'b001001_01010_01011_0000000000000000; // DIV  $11, $10
        memory[16] = 32'b000010_00000_01100_0000000000001001; // LW_3 $12, 9
        memory[17] = 32'b000010_00000_01101_0000000000001001; // LW_3 $13, 9
        memory[18] = 32'b001010_01100_01101_0000000000000000; // AND  $13, $12
        memory[19] = 32'b000010_00000_01110_0000000000010101; // LW_3 $14, 21
        memory[20] = 32'b000010_00000_01111_0000000000010010; // LW_3 $15, 18
        memory[21] = 32'b001011_01110_01111_0000000000010111; // OR   $15, $14
        memory[22] = 32'b000010_00000_10000_0000000000000011; // LW_3 $16, 3
        memory[23] = 32'b000010_00000_10001_0000000000000010; // LW_3 $17, 2
        memory[24] = 32'b001100_10001_10000_0000000000000000; // SHL   $16, $17
        memory[25] = 32'b000010_00000_10010_0000000000011000; // LW_3 $18, 24
        memory[26] = 32'b000010_00000_10011_0000000000000011; // LW_3 $19, 3
        memory[27] = 32'b001101_10011_10010_0000000000000000; // SHR   $18, $19
        memory[28] = 32'b000010_00000_10100_1111111111111000; // LW_3 $20, 65528
        memory[29] = 32'b001111_00000_10100_0000000000000000; // NOT  $20
        memory[30] = 32'b000010_00000_10101_0000000000101001; // LW_3 $21, 41
        memory[31] = 32'b010000_10101_00000_0000000000000000; // JR  $21
        memory[41] = 32'b010001_00000_00000_0000000000000101; // JPC PC + 5
        memory[47] = 32'b000010_00000_10110_0000000001100100; // LW_3 $22, 100
        memory[48] = 32'b010011_10110_00000_0000000000000000; // CALL ($22)
        memory[100] = 32'b001000_01000_01001_0000000000000000; // MUL  $9, $8
        memory[101] = 32'b010100_00000_00000_0000000000000000; // RET
        memory[49] = 32'b000010_00000_10111_0111111111111111; // LW_3 $23, 32767
        memory[50] = 32'b001000_10111_10111_0000000000000000; // MUL  $23, $23
        memory[51] = 32'b001000_10111_10111_0000000000000000; // MUL  $23, $23
        memory[52] = 32'b001000_10001_10111_0000000000000000; // MUL  $23, $17
        memory[53] = 32'b000010_00000_11000_0000000000000101; // LW_3 $24, 5
        memory[54] = 32'b000001_11000_11001_0000000000000000; // LW_2 $25, ($24)
        memory[55] = 32'b000110_11001_11001_0000000000000000; // ADD  $25, $25
        memory[56] = 32'b000010_00000_11000_0000000000000110; // LW_3 $24, 6
        memory[57] = 32'b000001_11000_11001_0000000000000000; // LW_2 $25, ($24)
        memory[58] = 32'b000010_00000_11000_0000000000000001; // LW_3 $24, 1
        memory[59] = 32'b000111_11001_11000_0000000000000000; // SUB  $24, $25
        memory[60] = 32'b000010_00000_11000_0000000000000100; // LW_3 $24, 4
        memory[61] = 32'b000001_11000_11001_0000000000000000; // LW_2 $25, ($24)
        memory[62] = 32'b001001_11001_11010_0000000000000000; // DIV  $26, $25
        memory[63] = 32'b000010_00000_11001_0000000000000100; // LW_3 $25, 4
        memory[64] = 32'b001110_11000_11001_0000000000000100; // CMP  $25, $24
        memory[65] = 32'b000010_00000_11001_0000000000000011; // LW_3 $25, 3
        memory[66] = 32'b001110_11000_11001_0000000000000100; // CMP  $25, $24
        memory[67] = 32'b000010_00000_11000_0000000000000010; // LW_3 $24, 2
        memory[68] = 32'b010101_00000_00000_0000000000000000; // NOP
        memory[69] = 32'b000010_00000_11010_0000000001100110; // LW_3 $26, 102
        memory[70] = 32'b001110_11000_11001_0000000000000100; // CMP  $25, $24        
        memory[71] = 32'b010010_11010_00000_0000000010000100; // BRFL ($26),00100
        memory[102] = 32'b010101_00000_00000_0000000000000000; // NOP
        memory[103] = 32'b000010_00000_11010_0000000001111000; // LW_3 $26, 120
        memory[104] = 32'b010011_11010_00000_0000000000000000; // CALL ($26)
        memory[120] = 32'b000010_00000_11010_0000000010010110; // LW_3 $26, 150
        memory[121] = 32'b010011_11010_00000_0000000000000000; // CALL ($26)
        memory[150] = 32'b000010_00000_11010_0000000011001000; // LW_3 $26, 200
        memory[151] = 32'b010011_11010_00000_0000000000000000; // CALL ($26)
        memory[200] = 32'b010101_00000_00000_0000000000000000; // NOP
        memory[201] = 32'b010100_00000_00000_0000000000000000; // RET
        memory[152] = 32'b010101_00000_00000_0000000000000000; // NOP
        memory[153] = 32'b010100_00000_00000_0000000000000000; // RET
        memory[122] = 32'b010101_00000_00000_0000000000000000; // NOP 
        memory[123] = 32'b010100_00000_00000_0000000000000000; // RET
        memory[105] = 32'b010101_00000_00000_0000000000000000; // NOP 
        // Adicione outras instrucoes aqui conforme necessario
    end

    always @ (posedge clk) begin
        instruction <= memory[address];
    end

endmodule
