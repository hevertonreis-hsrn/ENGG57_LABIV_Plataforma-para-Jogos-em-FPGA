module ControleInterface(
	input clock,
	input reset_n,
	input write,
	input read,
	input [31:0] writedata,
	output [31:0] readdata,
);

endmodule