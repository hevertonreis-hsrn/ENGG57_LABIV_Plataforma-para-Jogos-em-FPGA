	component EmbarcadoVGA is
		port (
			clk_clk                   : in    std_logic                     := 'X';             -- clk
			master_conduit_fifo_full  : in    std_logic                     := 'X';             -- fifo_full
			master_conduit_fifo_wr_en : out   std_logic;                                        -- fifo_wr_en
			master_conduit_exportdata : out   std_logic_vector(15 downto 0);                    -- exportdata
			master_conduit_pll_locked : in    std_logic                     := 'X';             -- pll_locked
			master_conduit_fifo_used  : in    std_logic_vector(8 downto 0)  := (others => 'X'); -- fifo_used
			master_conduit_fifo_empty : in    std_logic                     := 'X';             -- fifo_empty
			reset_reset_n             : in    std_logic                     := 'X';             -- reset_n
			sdram_addr                : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_ba                  : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_cas_n               : out   std_logic;                                        -- cas_n
			sdram_cke                 : out   std_logic;                                        -- cke
			sdram_cs_n                : out   std_logic;                                        -- cs_n
			sdram_dq                  : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_dqm                 : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_ras_n               : out   std_logic;                                        -- ras_n
			sdram_we_n                : out   std_logic;                                        -- we_n
			sw_conduit_export         : in    std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component EmbarcadoVGA;

	u0 : component EmbarcadoVGA
		port map (
			clk_clk                   => CONNECTED_TO_clk_clk,                   --            clk.clk
			master_conduit_fifo_full  => CONNECTED_TO_master_conduit_fifo_full,  -- master_conduit.fifo_full
			master_conduit_fifo_wr_en => CONNECTED_TO_master_conduit_fifo_wr_en, --               .fifo_wr_en
			master_conduit_exportdata => CONNECTED_TO_master_conduit_exportdata, --               .exportdata
			master_conduit_pll_locked => CONNECTED_TO_master_conduit_pll_locked, --               .pll_locked
			master_conduit_fifo_used  => CONNECTED_TO_master_conduit_fifo_used,  --               .fifo_used
			master_conduit_fifo_empty => CONNECTED_TO_master_conduit_fifo_empty, --               .fifo_empty
			reset_reset_n             => CONNECTED_TO_reset_reset_n,             --          reset.reset_n
			sdram_addr                => CONNECTED_TO_sdram_addr,                --          sdram.addr
			sdram_ba                  => CONNECTED_TO_sdram_ba,                  --               .ba
			sdram_cas_n               => CONNECTED_TO_sdram_cas_n,               --               .cas_n
			sdram_cke                 => CONNECTED_TO_sdram_cke,                 --               .cke
			sdram_cs_n                => CONNECTED_TO_sdram_cs_n,                --               .cs_n
			sdram_dq                  => CONNECTED_TO_sdram_dq,                  --               .dq
			sdram_dqm                 => CONNECTED_TO_sdram_dqm,                 --               .dqm
			sdram_ras_n               => CONNECTED_TO_sdram_ras_n,               --               .ras_n
			sdram_we_n                => CONNECTED_TO_sdram_we_n,                --               .we_n
			sw_conduit_export         => CONNECTED_TO_sw_conduit_export          --     sw_conduit.export
		);

