// EmbarcadoVGA_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module EmbarcadoVGA_tb (
	);

	wire         embarcadovga_inst_clk_bfm_clk_clk;       // EmbarcadoVGA_inst_clk_bfm:clk -> [EmbarcadoVGA_inst:clk_clk, EmbarcadoVGA_inst_reset_bfm:clk, sdram_controller_my_partner:clk]
	wire         embarcadovga_inst_sdram_cs_n;            // EmbarcadoVGA_inst:sdram_cs_n -> sdram_controller_my_partner:zs_cs_n
	wire   [3:0] embarcadovga_inst_sdram_dqm;             // EmbarcadoVGA_inst:sdram_dqm -> sdram_controller_my_partner:zs_dqm
	wire         embarcadovga_inst_sdram_cas_n;           // EmbarcadoVGA_inst:sdram_cas_n -> sdram_controller_my_partner:zs_cas_n
	wire         embarcadovga_inst_sdram_ras_n;           // EmbarcadoVGA_inst:sdram_ras_n -> sdram_controller_my_partner:zs_ras_n
	wire         embarcadovga_inst_sdram_we_n;            // EmbarcadoVGA_inst:sdram_we_n -> sdram_controller_my_partner:zs_we_n
	wire  [12:0] embarcadovga_inst_sdram_addr;            // EmbarcadoVGA_inst:sdram_addr -> sdram_controller_my_partner:zs_addr
	wire         embarcadovga_inst_sdram_cke;             // EmbarcadoVGA_inst:sdram_cke -> sdram_controller_my_partner:zs_cke
	wire  [31:0] embarcadovga_inst_sdram_dq;              // [] -> [EmbarcadoVGA_inst:sdram_dq, sdram_controller_my_partner:zs_dq]
	wire   [1:0] embarcadovga_inst_sdram_ba;              // EmbarcadoVGA_inst:sdram_ba -> sdram_controller_my_partner:zs_ba
	wire         embarcadovga_inst_reset_bfm_reset_reset; // EmbarcadoVGA_inst_reset_bfm:reset -> EmbarcadoVGA_inst:reset_reset_n

	EmbarcadoVGA embarcadovga_inst (
		.clk_clk       (embarcadovga_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (embarcadovga_inst_reset_bfm_reset_reset), // reset.reset_n
		.sdram_addr    (embarcadovga_inst_sdram_addr),            // sdram.addr
		.sdram_ba      (embarcadovga_inst_sdram_ba),              //      .ba
		.sdram_cas_n   (embarcadovga_inst_sdram_cas_n),           //      .cas_n
		.sdram_cke     (embarcadovga_inst_sdram_cke),             //      .cke
		.sdram_cs_n    (embarcadovga_inst_sdram_cs_n),            //      .cs_n
		.sdram_dq      (embarcadovga_inst_sdram_dq),              //      .dq
		.sdram_dqm     (embarcadovga_inst_sdram_dqm),             //      .dqm
		.sdram_ras_n   (embarcadovga_inst_sdram_ras_n),           //      .ras_n
		.sdram_we_n    (embarcadovga_inst_sdram_we_n)             //      .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) embarcadovga_inst_clk_bfm (
		.clk (embarcadovga_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) embarcadovga_inst_reset_bfm (
		.reset (embarcadovga_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (embarcadovga_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_sdram_partner_module sdram_controller_my_partner (
		.clk      (embarcadovga_inst_clk_bfm_clk_clk), //     clk.clk
		.zs_dq    (embarcadovga_inst_sdram_dq),        // conduit.dq
		.zs_addr  (embarcadovga_inst_sdram_addr),      //        .addr
		.zs_ba    (embarcadovga_inst_sdram_ba),        //        .ba
		.zs_cas_n (embarcadovga_inst_sdram_cas_n),     //        .cas_n
		.zs_cke   (embarcadovga_inst_sdram_cke),       //        .cke
		.zs_cs_n  (embarcadovga_inst_sdram_cs_n),      //        .cs_n
		.zs_dqm   (embarcadovga_inst_sdram_dqm),       //        .dqm
		.zs_ras_n (embarcadovga_inst_sdram_ras_n),     //        .ras_n
		.zs_we_n  (embarcadovga_inst_sdram_we_n)       //        .we_n
	);

endmodule
