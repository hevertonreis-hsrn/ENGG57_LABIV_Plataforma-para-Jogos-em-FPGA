// EmbarcadoVGA.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module EmbarcadoVGA (
		input  wire        clk_clk,                     //              clk.clk
		input  wire        master_conduit_1_fifo_full,  // master_conduit_1.fifo_full
		output wire        master_conduit_1_fifo_wr_en, //                 .fifo_wr_en
		output wire [31:0] master_conduit_1_exportdata, //                 .exportdata
		input  wire        master_conduit_1_pll_locked, //                 .pll_locked
		input  wire        reset_reset_n,               //            reset.reset_n
		output wire [12:0] sdram_addr,                  //            sdram.addr
		output wire [1:0]  sdram_ba,                    //                 .ba
		output wire        sdram_cas_n,                 //                 .cas_n
		output wire        sdram_cke,                   //                 .cke
		output wire        sdram_cs_n,                  //                 .cs_n
		inout  wire [31:0] sdram_dq,                    //                 .dq
		output wire [3:0]  sdram_dqm,                   //                 .dqm
		output wire        sdram_ras_n,                 //                 .ras_n
		output wire        sdram_we_n                   //                 .we_n
	);

	wire         master_interface_avalon_chipselect;                  // master_interface:chipselect -> mm_interconnect_0:master_interface_avalon_chipselect
	wire         master_interface_avalon_waitrequest;                 // mm_interconnect_0:master_interface_avalon_waitrequest -> master_interface:waitrequest
	wire  [31:0] master_interface_avalon_readdata;                    // mm_interconnect_0:master_interface_avalon_readdata -> master_interface:readdata
	wire         master_interface_avalon_read;                        // master_interface:read -> mm_interconnect_0:master_interface_avalon_read
	wire   [3:0] master_interface_avalon_byteenable;                  // master_interface:byteenable -> mm_interconnect_0:master_interface_avalon_byteenable
	wire  [29:0] master_interface_avalon_address;                     // master_interface:address -> mm_interconnect_0:master_interface_avalon_address
	wire         master_interface_avalon_readdatavalid;               // mm_interconnect_0:master_interface_avalon_readdatavalid -> master_interface:readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;    // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_readdata;      // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;   // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_controller_s1_address;       // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;          // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_controller_s1_byteenable;    // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid; // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;         // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_controller_s1_writedata;     // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         rst_controller_reset_out_reset;                      // rst_controller:reset_out -> [master_interface:reset_n, mm_interconnect_0:master_interface_reset_reset_bridge_in_reset_reset, sdram_controller:reset_n]

	Master_Interface master_interface (
		.clk           (clk_clk),                               //   clock.clk
		.reset_n       (~rst_controller_reset_out_reset),       //   reset.reset_n
		.waitrequest   (master_interface_avalon_waitrequest),   //  avalon.waitrequest
		.readdatavalid (master_interface_avalon_readdatavalid), //        .readdatavalid
		.readdata      (master_interface_avalon_readdata),      //        .readdata
		.read          (master_interface_avalon_read),          //        .read
		.chipselect    (master_interface_avalon_chipselect),    //        .chipselect
		.byteenable    (master_interface_avalon_byteenable),    //        .byteenable
		.address       (master_interface_avalon_address),       //        .address
		.fifo_full     (master_conduit_1_fifo_full),            // conduit.fifo_full
		.fifo_wr_en    (master_conduit_1_fifo_wr_en),           //        .fifo_wr_en
		.exportdata    (master_conduit_1_exportdata),           //        .exportdata
		.pll_locked    (master_conduit_1_pll_locked)            //        .pll_locked
	);

	EmbarcadoVGA_sdram_controller sdram_controller (
		.clk            (clk_clk),                                             //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                     // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	EmbarcadoVGA_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                        (clk_clk),                                             //                                      clk_clk.clk
		.master_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // master_interface_reset_reset_bridge_in_reset.reset
		.master_interface_avalon_address                    (master_interface_avalon_address),                     //                      master_interface_avalon.address
		.master_interface_avalon_waitrequest                (master_interface_avalon_waitrequest),                 //                                             .waitrequest
		.master_interface_avalon_byteenable                 (master_interface_avalon_byteenable),                  //                                             .byteenable
		.master_interface_avalon_chipselect                 (master_interface_avalon_chipselect),                  //                                             .chipselect
		.master_interface_avalon_read                       (master_interface_avalon_read),                        //                                             .read
		.master_interface_avalon_readdata                   (master_interface_avalon_readdata),                    //                                             .readdata
		.master_interface_avalon_readdatavalid              (master_interface_avalon_readdatavalid),               //                                             .readdatavalid
		.sdram_controller_s1_address                        (mm_interconnect_0_sdram_controller_s1_address),       //                          sdram_controller_s1.address
		.sdram_controller_s1_write                          (mm_interconnect_0_sdram_controller_s1_write),         //                                             .write
		.sdram_controller_s1_read                           (mm_interconnect_0_sdram_controller_s1_read),          //                                             .read
		.sdram_controller_s1_readdata                       (mm_interconnect_0_sdram_controller_s1_readdata),      //                                             .readdata
		.sdram_controller_s1_writedata                      (mm_interconnect_0_sdram_controller_s1_writedata),     //                                             .writedata
		.sdram_controller_s1_byteenable                     (mm_interconnect_0_sdram_controller_s1_byteenable),    //                                             .byteenable
		.sdram_controller_s1_readdatavalid                  (mm_interconnect_0_sdram_controller_s1_readdatavalid), //                                             .readdatavalid
		.sdram_controller_s1_waitrequest                    (mm_interconnect_0_sdram_controller_s1_waitrequest),   //                                             .waitrequest
		.sdram_controller_s1_chipselect                     (mm_interconnect_0_sdram_controller_s1_chipselect)     //                                             .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
