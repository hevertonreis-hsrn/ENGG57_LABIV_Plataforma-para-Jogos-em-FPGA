// SistemaEmbarcado.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SistemaEmbarcado (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         processadorcentral_data_master_waitrequest;        // mm_interconnect_0:ProcessadorCentral_data_master_waitrequest -> ProcessadorCentral:d_waitrequest
	wire  [31:0] processadorcentral_data_master_readdata;           // mm_interconnect_0:ProcessadorCentral_data_master_readdata -> ProcessadorCentral:d_readdata
	wire         processadorcentral_data_master_read;               // ProcessadorCentral:d_read -> mm_interconnect_0:ProcessadorCentral_data_master_read
	wire  [31:0] processadorcentral_data_master_address;            // ProcessadorCentral:d_address -> mm_interconnect_0:ProcessadorCentral_data_master_address
	wire         processadorcentral_data_master_write;              // ProcessadorCentral:d_write -> mm_interconnect_0:ProcessadorCentral_data_master_write
	wire  [31:0] processadorcentral_data_master_writedata;          // ProcessadorCentral:d_writedata -> mm_interconnect_0:ProcessadorCentral_data_master_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;               // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                 // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire   [9:0] mm_interconnect_0_ram_s1_address;                  // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;               // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                    // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                    // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire  [31:0] processadorcentral_instruction_master_readdata;    // mm_interconnect_1:ProcessadorCentral_instruction_master_readdata -> ProcessadorCentral:i_readdata
	wire         processadorcentral_instruction_master_waitrequest; // mm_interconnect_1:ProcessadorCentral_instruction_master_waitrequest -> ProcessadorCentral:i_waitrequest
	wire  [31:0] processadorcentral_instruction_master_address;     // ProcessadorCentral:i_address -> mm_interconnect_1:ProcessadorCentral_instruction_master_address
	wire         processadorcentral_instruction_master_read;        // ProcessadorCentral:i_read -> mm_interconnect_1:ProcessadorCentral_instruction_master_read
	wire         mm_interconnect_1_rom_s1_chipselect;               // mm_interconnect_1:ROM_s1_chipselect -> ROM:chipselect
	wire  [31:0] mm_interconnect_1_rom_s1_readdata;                 // ROM:readdata -> mm_interconnect_1:ROM_s1_readdata
	wire         mm_interconnect_1_rom_s1_debugaccess;              // mm_interconnect_1:ROM_s1_debugaccess -> ROM:debugaccess
	wire   [9:0] mm_interconnect_1_rom_s1_address;                  // mm_interconnect_1:ROM_s1_address -> ROM:address
	wire   [3:0] mm_interconnect_1_rom_s1_byteenable;               // mm_interconnect_1:ROM_s1_byteenable -> ROM:byteenable
	wire         mm_interconnect_1_rom_s1_write;                    // mm_interconnect_1:ROM_s1_write -> ROM:write
	wire  [31:0] mm_interconnect_1_rom_s1_writedata;                // mm_interconnect_1:ROM_s1_writedata -> ROM:writedata
	wire         mm_interconnect_1_rom_s1_clken;                    // mm_interconnect_1:ROM_s1_clken -> ROM:clken
	wire         rst_controller_reset_out_reset;                    // rst_controller:reset_out -> [ProcessadorCentral:reset_n, RAM:reset, ROM:reset, mm_interconnect_0:ProcessadorCentral_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ProcessadorCentral_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                // rst_controller:reset_req -> [RAM:reset_req, ROM:reset_req, rst_translator:reset_req_in]

	CPU processadorcentral (
		.clk           (clk_clk),                                           //              clock.clk
		.reset_n       (~rst_controller_reset_out_reset),                   //              reset.reset_n
		.d_waitrequest (processadorcentral_data_master_waitrequest),        //        data_master.waitrequest
		.d_readdata    (processadorcentral_data_master_readdata),           //                   .readdata
		.d_read        (processadorcentral_data_master_read),               //                   .read
		.d_write       (processadorcentral_data_master_write),              //                   .write
		.d_address     (processadorcentral_data_master_address),            //                   .address
		.d_writedata   (processadorcentral_data_master_writedata),          //                   .writedata
		.i_address     (processadorcentral_instruction_master_address),     // instruction_master.address
		.i_read        (processadorcentral_instruction_master_read),        //                   .read
		.i_readdata    (processadorcentral_instruction_master_readdata),    //                   .readdata
		.i_waitrequest (processadorcentral_instruction_master_waitrequest)  //                   .waitrequest
	);

	SistemaEmbarcado_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	SistemaEmbarcado_ROM rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_1_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_1_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_1_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_1_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_1_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_1_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_1_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_1_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	SistemaEmbarcado_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                        (clk_clk),                                    //                                      clock_clk.clk
		.ProcessadorCentral_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),             // ProcessadorCentral_reset_reset_bridge_in_reset.reset
		.ProcessadorCentral_data_master_address               (processadorcentral_data_master_address),     //                 ProcessadorCentral_data_master.address
		.ProcessadorCentral_data_master_waitrequest           (processadorcentral_data_master_waitrequest), //                                               .waitrequest
		.ProcessadorCentral_data_master_read                  (processadorcentral_data_master_read),        //                                               .read
		.ProcessadorCentral_data_master_readdata              (processadorcentral_data_master_readdata),    //                                               .readdata
		.ProcessadorCentral_data_master_write                 (processadorcentral_data_master_write),       //                                               .write
		.ProcessadorCentral_data_master_writedata             (processadorcentral_data_master_writedata),   //                                               .writedata
		.RAM_s1_address                                       (mm_interconnect_0_ram_s1_address),           //                                         RAM_s1.address
		.RAM_s1_write                                         (mm_interconnect_0_ram_s1_write),             //                                               .write
		.RAM_s1_readdata                                      (mm_interconnect_0_ram_s1_readdata),          //                                               .readdata
		.RAM_s1_writedata                                     (mm_interconnect_0_ram_s1_writedata),         //                                               .writedata
		.RAM_s1_byteenable                                    (mm_interconnect_0_ram_s1_byteenable),        //                                               .byteenable
		.RAM_s1_chipselect                                    (mm_interconnect_0_ram_s1_chipselect),        //                                               .chipselect
		.RAM_s1_clken                                         (mm_interconnect_0_ram_s1_clken)              //                                               .clken
	);

	SistemaEmbarcado_mm_interconnect_1 mm_interconnect_1 (
		.clock_clk_clk                                        (clk_clk),                                           //                                      clock_clk.clk
		.ProcessadorCentral_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                    // ProcessadorCentral_reset_reset_bridge_in_reset.reset
		.ProcessadorCentral_instruction_master_address        (processadorcentral_instruction_master_address),     //          ProcessadorCentral_instruction_master.address
		.ProcessadorCentral_instruction_master_waitrequest    (processadorcentral_instruction_master_waitrequest), //                                               .waitrequest
		.ProcessadorCentral_instruction_master_read           (processadorcentral_instruction_master_read),        //                                               .read
		.ProcessadorCentral_instruction_master_readdata       (processadorcentral_instruction_master_readdata),    //                                               .readdata
		.ROM_s1_address                                       (mm_interconnect_1_rom_s1_address),                  //                                         ROM_s1.address
		.ROM_s1_write                                         (mm_interconnect_1_rom_s1_write),                    //                                               .write
		.ROM_s1_readdata                                      (mm_interconnect_1_rom_s1_readdata),                 //                                               .readdata
		.ROM_s1_writedata                                     (mm_interconnect_1_rom_s1_writedata),                //                                               .writedata
		.ROM_s1_byteenable                                    (mm_interconnect_1_rom_s1_byteenable),               //                                               .byteenable
		.ROM_s1_chipselect                                    (mm_interconnect_1_rom_s1_chipselect),               //                                               .chipselect
		.ROM_s1_clken                                         (mm_interconnect_1_rom_s1_clken),                    //                                               .clken
		.ROM_s1_debugaccess                                   (mm_interconnect_1_rom_s1_debugaccess)               //                                               .debugaccess
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
