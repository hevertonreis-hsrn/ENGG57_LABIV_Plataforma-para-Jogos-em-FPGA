// embedded_vpu_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module embedded_vpu_tb (
	);

	wire         embedded_vpu_inst_clk_bfm_clk_clk;                                  // embedded_vpu_inst_clk_bfm:clk -> [embedded_vpu_inst:clk_clk, embedded_vpu_inst_background_loader_conduit_bfm:clk, embedded_vpu_inst_composer_conduit_bfm:clk, embedded_vpu_inst_reset_bfm:clk, sdram_controller_my_partner:clk]
	wire   [0:0] embedded_vpu_inst_background_loader_conduit_bfm_conduit_pll_locked; // embedded_vpu_inst_background_loader_conduit_bfm:sig_pll_locked -> embedded_vpu_inst:background_loader_conduit_pll_locked
	wire         embedded_vpu_inst_composer_conduit_wrreq;                           // embedded_vpu_inst:composer_conduit_wrreq -> embedded_vpu_inst_composer_conduit_bfm:sig_wrreq
	wire  [23:0] embedded_vpu_inst_composer_conduit_pixel_out;                       // embedded_vpu_inst:composer_conduit_pixel_out -> embedded_vpu_inst_composer_conduit_bfm:sig_pixel_out
	wire   [0:0] embedded_vpu_inst_composer_conduit_bfm_conduit_wrfull;              // embedded_vpu_inst_composer_conduit_bfm:sig_wrfull -> embedded_vpu_inst:composer_conduit_wrfull
	wire   [3:0] embedded_vpu_inst_key_external_connection_bfm_conduit_export;       // embedded_vpu_inst_key_external_connection_bfm:sig_export -> embedded_vpu_inst:key_external_connection_export
	wire         embedded_vpu_inst_sdram_controller_wire_cs_n;                       // embedded_vpu_inst:sdram_controller_wire_cs_n -> sdram_controller_my_partner:zs_cs_n
	wire   [3:0] embedded_vpu_inst_sdram_controller_wire_dqm;                        // embedded_vpu_inst:sdram_controller_wire_dqm -> sdram_controller_my_partner:zs_dqm
	wire         embedded_vpu_inst_sdram_controller_wire_cas_n;                      // embedded_vpu_inst:sdram_controller_wire_cas_n -> sdram_controller_my_partner:zs_cas_n
	wire         embedded_vpu_inst_sdram_controller_wire_ras_n;                      // embedded_vpu_inst:sdram_controller_wire_ras_n -> sdram_controller_my_partner:zs_ras_n
	wire         embedded_vpu_inst_sdram_controller_wire_we_n;                       // embedded_vpu_inst:sdram_controller_wire_we_n -> sdram_controller_my_partner:zs_we_n
	wire  [12:0] embedded_vpu_inst_sdram_controller_wire_addr;                       // embedded_vpu_inst:sdram_controller_wire_addr -> sdram_controller_my_partner:zs_addr
	wire         embedded_vpu_inst_sdram_controller_wire_cke;                        // embedded_vpu_inst:sdram_controller_wire_cke -> sdram_controller_my_partner:zs_cke
	wire  [31:0] embedded_vpu_inst_sdram_controller_wire_dq;                         // [] -> [embedded_vpu_inst:sdram_controller_wire_dq, sdram_controller_my_partner:zs_dq]
	wire   [1:0] embedded_vpu_inst_sdram_controller_wire_ba;                         // embedded_vpu_inst:sdram_controller_wire_ba -> sdram_controller_my_partner:zs_ba
	wire         embedded_vpu_inst_reset_bfm_reset_reset;                            // embedded_vpu_inst_reset_bfm:reset -> [embedded_vpu_inst:reset_reset_n, embedded_vpu_inst_background_loader_conduit_bfm:reset, embedded_vpu_inst_composer_conduit_bfm:reset]

	embedded_vpu embedded_vpu_inst (
		.background_loader_conduit_pll_locked (embedded_vpu_inst_background_loader_conduit_bfm_conduit_pll_locked), // background_loader_conduit.pll_locked
		.clk_clk                              (embedded_vpu_inst_clk_bfm_clk_clk),                                  //                       clk.clk
		.composer_conduit_pixel_out           (embedded_vpu_inst_composer_conduit_pixel_out),                       //          composer_conduit.pixel_out
		.composer_conduit_wrfull              (embedded_vpu_inst_composer_conduit_bfm_conduit_wrfull),              //                          .wrfull
		.composer_conduit_wrreq               (embedded_vpu_inst_composer_conduit_wrreq),                           //                          .wrreq
		.key_external_connection_export       (embedded_vpu_inst_key_external_connection_bfm_conduit_export),       //   key_external_connection.export
		.reset_reset_n                        (embedded_vpu_inst_reset_bfm_reset_reset),                            //                     reset.reset_n
		.sdram_controller_wire_addr           (embedded_vpu_inst_sdram_controller_wire_addr),                       //     sdram_controller_wire.addr
		.sdram_controller_wire_ba             (embedded_vpu_inst_sdram_controller_wire_ba),                         //                          .ba
		.sdram_controller_wire_cas_n          (embedded_vpu_inst_sdram_controller_wire_cas_n),                      //                          .cas_n
		.sdram_controller_wire_cke            (embedded_vpu_inst_sdram_controller_wire_cke),                        //                          .cke
		.sdram_controller_wire_cs_n           (embedded_vpu_inst_sdram_controller_wire_cs_n),                       //                          .cs_n
		.sdram_controller_wire_dq             (embedded_vpu_inst_sdram_controller_wire_dq),                         //                          .dq
		.sdram_controller_wire_dqm            (embedded_vpu_inst_sdram_controller_wire_dqm),                        //                          .dqm
		.sdram_controller_wire_ras_n          (embedded_vpu_inst_sdram_controller_wire_ras_n),                      //                          .ras_n
		.sdram_controller_wire_we_n           (embedded_vpu_inst_sdram_controller_wire_we_n)                        //                          .we_n
	);

	altera_conduit_bfm embedded_vpu_inst_background_loader_conduit_bfm (
		.clk            (embedded_vpu_inst_clk_bfm_clk_clk),                                  //     clk.clk
		.reset          (~embedded_vpu_inst_reset_bfm_reset_reset),                           //   reset.reset
		.sig_pll_locked (embedded_vpu_inst_background_loader_conduit_bfm_conduit_pll_locked)  // conduit.pll_locked
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (100000000),
		.CLOCK_UNIT (1)
	) embedded_vpu_inst_clk_bfm (
		.clk (embedded_vpu_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0002 embedded_vpu_inst_composer_conduit_bfm (
		.clk           (embedded_vpu_inst_clk_bfm_clk_clk),                     //     clk.clk
		.reset         (~embedded_vpu_inst_reset_bfm_reset_reset),              //   reset.reset
		.sig_pixel_out (embedded_vpu_inst_composer_conduit_pixel_out),          // conduit.pixel_out
		.sig_wrfull    (embedded_vpu_inst_composer_conduit_bfm_conduit_wrfull), //        .wrfull
		.sig_wrreq     (embedded_vpu_inst_composer_conduit_wrreq)               //        .wrreq
	);

	altera_conduit_bfm_0003 embedded_vpu_inst_key_external_connection_bfm (
		.sig_export (embedded_vpu_inst_key_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) embedded_vpu_inst_reset_bfm (
		.reset (embedded_vpu_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (embedded_vpu_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_sdram_partner_module sdram_controller_my_partner (
		.clk      (embedded_vpu_inst_clk_bfm_clk_clk),             //     clk.clk
		.zs_dq    (embedded_vpu_inst_sdram_controller_wire_dq),    // conduit.dq
		.zs_addr  (embedded_vpu_inst_sdram_controller_wire_addr),  //        .addr
		.zs_ba    (embedded_vpu_inst_sdram_controller_wire_ba),    //        .ba
		.zs_cas_n (embedded_vpu_inst_sdram_controller_wire_cas_n), //        .cas_n
		.zs_cke   (embedded_vpu_inst_sdram_controller_wire_cke),   //        .cke
		.zs_cs_n  (embedded_vpu_inst_sdram_controller_wire_cs_n),  //        .cs_n
		.zs_dqm   (embedded_vpu_inst_sdram_controller_wire_dqm),   //        .dqm
		.zs_ras_n (embedded_vpu_inst_sdram_controller_wire_ras_n), //        .ras_n
		.zs_we_n  (embedded_vpu_inst_sdram_controller_wire_we_n)   //        .we_n
	);

endmodule
