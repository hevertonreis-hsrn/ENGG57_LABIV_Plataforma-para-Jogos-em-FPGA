// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Sat Apr 19 16:35:05 2025"

module ModuloProcessador(
	clk,
	rst
);


input wire	clk;
input wire	rst;

wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	[7:0] SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_62;
wire	[4:0] SYNTHESIZED_WIRE_63;
wire	[4:0] SYNTHESIZED_WIRE_9;
wire	[4:0] SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_14;
wire	[31:0] SYNTHESIZED_WIRE_15;
wire	[7:0] SYNTHESIZED_WIRE_16;
wire	[31:0] SYNTHESIZED_WIRE_65;
wire	[4:0] SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	[31:0] SYNTHESIZED_WIRE_66;
wire	[1:0] SYNTHESIZED_WIRE_28;
wire	[1:0] SYNTHESIZED_WIRE_29;
wire	[5:0] SYNTHESIZED_WIRE_30;
wire	[7:0] SYNTHESIZED_WIRE_31;
wire	[31:0] SYNTHESIZED_WIRE_32;
wire	[31:0] SYNTHESIZED_WIRE_33;
wire	[31:0] SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_67;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	[31:0] SYNTHESIZED_WIRE_44;
wire	[4:0] SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	[31:0] SYNTHESIZED_WIRE_48;
wire	[31:0] SYNTHESIZED_WIRE_49;
wire	[4:0] SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_52;
wire	[4:0] SYNTHESIZED_WIRE_56;





IF_STAGE	b2v_inst(
	.clk_Mem(clk),
	.clk(SYNTHESIZED_WIRE_59),
	.rst(SYNTHESIZED_WIRE_60),
	.PCSrc(SYNTHESIZED_WIRE_61),
	.HD_HoldPC(SYNTHESIZED_WIRE_3),
	.HD_Hold_IF_ID(SYNTHESIZED_WIRE_4),
	.IF_Flush(SYNTHESIZED_WIRE_61),
	.BranchTarget(SYNTHESIZED_WIRE_6),
	.IF_ID_Inst(SYNTHESIZED_WIRE_15),
	.IF_ID_PC(SYNTHESIZED_WIRE_16));


HazardDetectionUnit	b2v_inst1(
	.ID_EX_MemRead(SYNTHESIZED_WIRE_62),
	.ID_EX_WriteReg(SYNTHESIZED_WIRE_63),
	.r1(SYNTHESIZED_WIRE_9),
	.r2(SYNTHESIZED_WIRE_10),
	.HD_HoldPC(SYNTHESIZED_WIRE_3),
	.HD_Hold_IF_ID(SYNTHESIZED_WIRE_4),
	.HD_HoldControl(SYNTHESIZED_WIRE_14));


ID_STAGE	b2v_inst2(
	.clk(SYNTHESIZED_WIRE_59),
	.rst(SYNTHESIZED_WIRE_60),
	.RegWrite(SYNTHESIZED_WIRE_64),
	.clk_Mem(clk),
	.HD_HoldControl(SYNTHESIZED_WIRE_14),
	.IF_ID_Inst(SYNTHESIZED_WIRE_15),
	.IF_ID_PC(SYNTHESIZED_WIRE_16),
	.WriteData(SYNTHESIZED_WIRE_65),
	.WriteReg(SYNTHESIZED_WIRE_18),
	.ID_EX_MemToReg(SYNTHESIZED_WIRE_21),
	.ID_EX_RegWrite(SYNTHESIZED_WIRE_22),
	.ID_EX_Branch(SYNTHESIZED_WIRE_23),
	.ID_EX_MemRead(SYNTHESIZED_WIRE_62),
	.ID_EX_MemWrite(SYNTHESIZED_WIRE_25),
	.ID_EX_ALUSrc(SYNTHESIZED_WIRE_26),
	.ID_EX_ALUOp(SYNTHESIZED_WIRE_30),
	.ID_EX_BranchTarget(SYNTHESIZED_WIRE_31),
	.ID_EX_ReadData1(SYNTHESIZED_WIRE_32),
	.ID_EX_ReadData2(SYNTHESIZED_WIRE_33),
	.ID_EX_Rs(SYNTHESIZED_WIRE_56),
	.ID_EX_SignExtImm(SYNTHESIZED_WIRE_34),
	.ID_EX_WriteReg(SYNTHESIZED_WIRE_63),
	.r1(SYNTHESIZED_WIRE_9),
	.r2(SYNTHESIZED_WIRE_10));


EX_STAGE	b2v_inst3(
	.clk(SYNTHESIZED_WIRE_59),
	.rst(SYNTHESIZED_WIRE_60),
	.ID_EX_MemToReg(SYNTHESIZED_WIRE_21),
	.ID_EX_RegWrite(SYNTHESIZED_WIRE_22),
	.ID_EX_Branch(SYNTHESIZED_WIRE_23),
	.ID_EX_MemRead(SYNTHESIZED_WIRE_62),
	.ID_EX_MemWrite(SYNTHESIZED_WIRE_25),
	.ID_EX_ALUSrc(SYNTHESIZED_WIRE_26),
	.EX_Data(SYNTHESIZED_WIRE_66),
	.FowardA(SYNTHESIZED_WIRE_28),
	.FowardB(SYNTHESIZED_WIRE_29),
	.ID_EX_ALUOp(SYNTHESIZED_WIRE_30),
	.ID_EX_BranchTarget(SYNTHESIZED_WIRE_31),
	.ID_EX_ReadData1(SYNTHESIZED_WIRE_32),
	.ID_EX_ReadData2(SYNTHESIZED_WIRE_33),
	.ID_EX_SignExtImm(SYNTHESIZED_WIRE_34),
	.ID_EX_WriteReg(SYNTHESIZED_WIRE_63),
	.MEM_Data(SYNTHESIZED_WIRE_65),
	.BranchTaken(SYNTHESIZED_WIRE_61),
	.EX_MEM_MemToReg(SYNTHESIZED_WIRE_39),
	.EX_MEM_RegWrite(SYNTHESIZED_WIRE_67),
	.EX_MEM_MemRead(SYNTHESIZED_WIRE_41),
	.EX_MEM_MemWrite(SYNTHESIZED_WIRE_42),
	.BranchTarget(SYNTHESIZED_WIRE_6),
	.EX_MEM_ALUResult(SYNTHESIZED_WIRE_66),
	.EX_MEM_WriteData(SYNTHESIZED_WIRE_44),
	.EX_MEM_WriteReg(SYNTHESIZED_WIRE_68));


MEM_STAGE	b2v_inst4(
	.clk_Mem(clk),
	.clk(SYNTHESIZED_WIRE_59),
	.rst(SYNTHESIZED_WIRE_60),
	.EX_MEM_MemToReg(SYNTHESIZED_WIRE_39),
	.EX_MEM_RegWrite(SYNTHESIZED_WIRE_67),
	.EX_MEM_MemRead(SYNTHESIZED_WIRE_41),
	.EX_MEM_MemWrite(SYNTHESIZED_WIRE_42),
	.EX_MEM_ALUResult(SYNTHESIZED_WIRE_66),
	.EX_MEM_WriteData(SYNTHESIZED_WIRE_44),
	.EX_MEM_WriteReg(SYNTHESIZED_WIRE_68),
	.MEM_WB_RegWrite(SYNTHESIZED_WIRE_46),
	.MEM_WB_MemToReg(SYNTHESIZED_WIRE_47),
	.MEM_WB_ALUResult(SYNTHESIZED_WIRE_48),
	.MEM_WB_ReadData(SYNTHESIZED_WIRE_49),
	.MEM_WB_WriteReg(SYNTHESIZED_WIRE_69));


WB_STAGE	b2v_inst5(
	.MEM_WB_RegWrite(SYNTHESIZED_WIRE_46),
	.MEM_WB_MemToReg(SYNTHESIZED_WIRE_47),
	.MEM_WB_ALUResult(SYNTHESIZED_WIRE_48),
	.MEM_WB_ReadData(SYNTHESIZED_WIRE_49),
	.MEM_WB_WriteReg(SYNTHESIZED_WIRE_69),
	.RegWrite(SYNTHESIZED_WIRE_64),
	.WriteData(SYNTHESIZED_WIRE_65),
	.WriteReg(SYNTHESIZED_WIRE_18));


DividerPLL	b2v_inst6(
	.inclk0(clk),
	.areset(rst),
	.c0(SYNTHESIZED_WIRE_59));


ResetSync	b2v_inst7(
	.clk(SYNTHESIZED_WIRE_59),
	.rst_async(SYNTHESIZED_WIRE_52),
	.rst_sync(SYNTHESIZED_WIRE_60));


ForwardingUnit	b2v_inst8(
	.EX_MEM_RegWrite(SYNTHESIZED_WIRE_67),
	.MEM_WB_RegWrite(SYNTHESIZED_WIRE_64),
	.EX_MEM_rd(SYNTHESIZED_WIRE_68),
	.ID_EX_rs1(SYNTHESIZED_WIRE_56),
	.ID_EX_rs2(SYNTHESIZED_WIRE_63),
	.MEM_WB_rd(SYNTHESIZED_WIRE_69),
	.ForwardA(SYNTHESIZED_WIRE_28),
	.ForwardB(SYNTHESIZED_WIRE_29));

assign	SYNTHESIZED_WIRE_52 =  ~rst;


endmodule
