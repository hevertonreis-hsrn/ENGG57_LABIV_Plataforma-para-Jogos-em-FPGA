// EmbarcadoVGA_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module EmbarcadoVGA_tb (
	);

	wire         embarcadovga_inst_clk_bfm_clk_clk;                       // EmbarcadoVGA_inst_clk_bfm:clk -> [EmbarcadoVGA_inst:clk_clk, EmbarcadoVGA_inst_master_conduit_bfm:clk, EmbarcadoVGA_inst_reset_bfm:clk, sdram_controller_my_partner:clk]
	wire  [15:0] embarcadovga_inst_master_conduit_exportdata;             // EmbarcadoVGA_inst:master_conduit_exportdata -> EmbarcadoVGA_inst_master_conduit_bfm:sig_exportdata
	wire   [0:0] embarcadovga_inst_master_conduit_bfm_conduit_fifo_full;  // EmbarcadoVGA_inst_master_conduit_bfm:sig_fifo_full -> EmbarcadoVGA_inst:master_conduit_fifo_full
	wire         embarcadovga_inst_master_conduit_fifo_wr_en;             // EmbarcadoVGA_inst:master_conduit_fifo_wr_en -> EmbarcadoVGA_inst_master_conduit_bfm:sig_fifo_wr_en
	wire   [0:0] embarcadovga_inst_master_conduit_bfm_conduit_fifo_empty; // EmbarcadoVGA_inst_master_conduit_bfm:sig_fifo_empty -> EmbarcadoVGA_inst:master_conduit_fifo_empty
	wire   [8:0] embarcadovga_inst_master_conduit_bfm_conduit_fifo_used;  // EmbarcadoVGA_inst_master_conduit_bfm:sig_fifo_used -> EmbarcadoVGA_inst:master_conduit_fifo_used
	wire   [0:0] embarcadovga_inst_master_conduit_bfm_conduit_pll_locked; // EmbarcadoVGA_inst_master_conduit_bfm:sig_pll_locked -> EmbarcadoVGA_inst:master_conduit_pll_locked
	wire         embarcadovga_inst_sdram_cs_n;                            // EmbarcadoVGA_inst:sdram_cs_n -> sdram_controller_my_partner:zs_cs_n
	wire   [1:0] embarcadovga_inst_sdram_dqm;                             // EmbarcadoVGA_inst:sdram_dqm -> sdram_controller_my_partner:zs_dqm
	wire         embarcadovga_inst_sdram_cas_n;                           // EmbarcadoVGA_inst:sdram_cas_n -> sdram_controller_my_partner:zs_cas_n
	wire         embarcadovga_inst_sdram_ras_n;                           // EmbarcadoVGA_inst:sdram_ras_n -> sdram_controller_my_partner:zs_ras_n
	wire         embarcadovga_inst_sdram_we_n;                            // EmbarcadoVGA_inst:sdram_we_n -> sdram_controller_my_partner:zs_we_n
	wire  [12:0] embarcadovga_inst_sdram_addr;                            // EmbarcadoVGA_inst:sdram_addr -> sdram_controller_my_partner:zs_addr
	wire         embarcadovga_inst_sdram_cke;                             // EmbarcadoVGA_inst:sdram_cke -> sdram_controller_my_partner:zs_cke
	wire  [15:0] embarcadovga_inst_sdram_dq;                              // [] -> [EmbarcadoVGA_inst:sdram_dq, sdram_controller_my_partner:zs_dq]
	wire   [1:0] embarcadovga_inst_sdram_ba;                              // EmbarcadoVGA_inst:sdram_ba -> sdram_controller_my_partner:zs_ba
	wire   [1:0] embarcadovga_inst_sw_conduit_bfm_conduit_export;         // EmbarcadoVGA_inst_sw_conduit_bfm:sig_export -> EmbarcadoVGA_inst:sw_conduit_export
	wire         embarcadovga_inst_reset_bfm_reset_reset;                 // EmbarcadoVGA_inst_reset_bfm:reset -> [EmbarcadoVGA_inst:reset_reset_n, EmbarcadoVGA_inst_master_conduit_bfm:reset]

	EmbarcadoVGA embarcadovga_inst (
		.clk_clk                   (embarcadovga_inst_clk_bfm_clk_clk),                       //            clk.clk
		.master_conduit_fifo_full  (embarcadovga_inst_master_conduit_bfm_conduit_fifo_full),  // master_conduit.fifo_full
		.master_conduit_fifo_wr_en (embarcadovga_inst_master_conduit_fifo_wr_en),             //               .fifo_wr_en
		.master_conduit_exportdata (embarcadovga_inst_master_conduit_exportdata),             //               .exportdata
		.master_conduit_pll_locked (embarcadovga_inst_master_conduit_bfm_conduit_pll_locked), //               .pll_locked
		.master_conduit_fifo_used  (embarcadovga_inst_master_conduit_bfm_conduit_fifo_used),  //               .fifo_used
		.master_conduit_fifo_empty (embarcadovga_inst_master_conduit_bfm_conduit_fifo_empty), //               .fifo_empty
		.reset_reset_n             (embarcadovga_inst_reset_bfm_reset_reset),                 //          reset.reset_n
		.sdram_addr                (embarcadovga_inst_sdram_addr),                            //          sdram.addr
		.sdram_ba                  (embarcadovga_inst_sdram_ba),                              //               .ba
		.sdram_cas_n               (embarcadovga_inst_sdram_cas_n),                           //               .cas_n
		.sdram_cke                 (embarcadovga_inst_sdram_cke),                             //               .cke
		.sdram_cs_n                (embarcadovga_inst_sdram_cs_n),                            //               .cs_n
		.sdram_dq                  (embarcadovga_inst_sdram_dq),                              //               .dq
		.sdram_dqm                 (embarcadovga_inst_sdram_dqm),                             //               .dqm
		.sdram_ras_n               (embarcadovga_inst_sdram_ras_n),                           //               .ras_n
		.sdram_we_n                (embarcadovga_inst_sdram_we_n),                            //               .we_n
		.sw_conduit_export         (embarcadovga_inst_sw_conduit_bfm_conduit_export)          //     sw_conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (100000000),
		.CLOCK_UNIT (1)
	) embarcadovga_inst_clk_bfm (
		.clk (embarcadovga_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm embarcadovga_inst_master_conduit_bfm (
		.clk            (embarcadovga_inst_clk_bfm_clk_clk),                       //     clk.clk
		.reset          (~embarcadovga_inst_reset_bfm_reset_reset),                //   reset.reset
		.sig_exportdata (embarcadovga_inst_master_conduit_exportdata),             // conduit.exportdata
		.sig_fifo_empty (embarcadovga_inst_master_conduit_bfm_conduit_fifo_empty), //        .fifo_empty
		.sig_fifo_full  (embarcadovga_inst_master_conduit_bfm_conduit_fifo_full),  //        .fifo_full
		.sig_fifo_used  (embarcadovga_inst_master_conduit_bfm_conduit_fifo_used),  //        .fifo_used
		.sig_fifo_wr_en (embarcadovga_inst_master_conduit_fifo_wr_en),             //        .fifo_wr_en
		.sig_pll_locked (embarcadovga_inst_master_conduit_bfm_conduit_pll_locked)  //        .pll_locked
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) embarcadovga_inst_reset_bfm (
		.reset (embarcadovga_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (embarcadovga_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0002 embarcadovga_inst_sw_conduit_bfm (
		.sig_export (embarcadovga_inst_sw_conduit_bfm_conduit_export)  // conduit.export
	);

	altera_sdram_partner_module sdram_controller_my_partner (
		.clk      (embarcadovga_inst_clk_bfm_clk_clk), //     clk.clk
		.zs_dq    (embarcadovga_inst_sdram_dq),        // conduit.dq
		.zs_addr  (embarcadovga_inst_sdram_addr),      //        .addr
		.zs_ba    (embarcadovga_inst_sdram_ba),        //        .ba
		.zs_cas_n (embarcadovga_inst_sdram_cas_n),     //        .cas_n
		.zs_cke   (embarcadovga_inst_sdram_cke),       //        .cke
		.zs_cs_n  (embarcadovga_inst_sdram_cs_n),      //        .cs_n
		.zs_dqm   (embarcadovga_inst_sdram_dqm),       //        .dqm
		.zs_ras_n (embarcadovga_inst_sdram_ras_n),     //        .ras_n
		.zs_we_n  (embarcadovga_inst_sdram_we_n)       //        .we_n
	);

endmodule
